//Verilog HDL for "VIS015libraryRAW", "ARD00timerclockRAW1" "functional"


module ARD00timerclockRAW1 ( C0, C1, tdo_timerclock, timerclock, G, V, en, ten_timerclock
);

  input V;
  output timerclock;
  output tdo_timerclock;
  input ten_timerclock;
  input en;
  input G;
  output C1;
  output C0;
endmodule
