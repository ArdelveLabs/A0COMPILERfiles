//Verilog HDL for "VIS015libraryRAW", "ARD00referenceRAW2" "functional"


module ARD00referenceRAW2 ( V, G, R, trimREF );

  input  [4:0] trimREF;
  input V;
  inout  [5:0] R;
  input G;
endmodule
