//Verilog HDL for "VIS015libraryRAW", "ARD00timerclockRAW2" "functional"


module ARD00timerclockRAW2 ( V, CN0, CN1, CN2, CN3, trimTIMERCLOCK, G );

  input CN0;
  input V;
  input CN1;
  input  [3:0] trimTIMERCLOCK;
  input CN2;
  input G;
  input CN3;
endmodule
